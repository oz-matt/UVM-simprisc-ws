	
package instruction_sequences;
	
	`include "src/seq_items/instruction_base_si.sv"
	`include "src/seq_items/arithmetic_instruction_si.sv"
	`include "src/seq_items/store_instruction_si.sv"
	`include "src/seq_items/load_instruction_si.sv"
	
endpackage