`ifndef RISCV_INSTRUCTION_PROPERTIES
`define RISCV_INSTRUCTION_PROPERTIES

package riscv_instruction_properties;
	
	typedef enum bit [4:0] {
		RV32I,
		RV64I,
		RV32M,
		RV64M,
		RV32A,
		RV64A,
		RV32F,
		RV32FC,
		RV64F,
		RV32D,
		RV32DC,
		RV64D,
		RV32C,
		RV64C,
		RV128I,
		RV128C
	} riscv_instr_group_t;

	typedef enum {
		// RV32I instructions
		LUI,
		AUIPC,
		JAL,
		JALR,
		BEQ,
		BNE,
		BLT,
		BGE,
		BLTU,
		BGEU,
		LB,
		LH,
		LW,
		LBU,
		LHU,
		SB,
		SH,
		SW,
		ADDI,
		SLTI,
		SLTIU,
		XORI,
		ORI,
		ANDI,
		SLLI,
		SRLI,
		SRAI,
		ADD,
		SUB,
		SLL,
		SLT,
		SLTU,
		XOR,
		SRL,
		SRA,
		OR,
		AND,
		NOP,
		FENCE,
		FENCEI,
		ECALL,
		EBREAK,
		CSRRW,
		CSRRS,
		CSRRC,
		CSRRWI,
		CSRRSI,
		CSRRCI,
		// RV32M instructions
		MUL,
		MULH,
		MULHSU,
		MULHU,
		DIV,
		DIVU,
		REM,
		REMU,
		// RV64M instructions
		MULW,
		DIVW,
		DIVUW,
		REMW,
		REMUW,
		// RV32F instructions
		FLW,
		FSW,
		FMADD_S,
		FMSUB_S,
		FNMSUB_S,
		FNMADD_S,
		FADD_S,
		FSUB_S,
		FMUL_S,
		FDIV_S,
		FSQRT_S,
		FSGNJ_S,
		FSGNJN_S,
		FSGNJX_S,
		FMIN_S,
		FMAX_S,
		FCVT_W_S,
		FCVT_WU_S,
		FMV_X_W,
		FEQ_S,
		FLT_S,
		FLE_S,
		FCLASS_S,
		FCVT_S_W,
		FCVT_S_WU,
		FMV_W_X,
		FCVT_L_S,
		FCVT_LU_S,
		FCVT_S_L,
		FCVT_S_LU,
		// RV64I
		LWU,
		LD,
		SD,
		ADDIW,
		SLLIW,
		SRLIW,
		SRAIW,
		ADDW,
		SUBW,
		SLLW,
		SRLW,
		SRAW,
		// RV32C
		C_LW,
		C_SW,
		C_LWSP,
		C_SWSP,
		C_ADDI4SPN,
		C_ADDI,
		C_LI,
		C_ADDI16SP,
		C_LUI,
		C_SRLI,
		C_SRAI,
		C_ANDI,
		C_SUB,
		C_XOR,
		C_OR,
		C_AND,
		C_BEQZ,
		C_BNEZ,
		C_SLLI,
		C_MV,
		C_EBREAK,
		C_ADD,
		C_NOP,
		C_J,
		C_JAL,
		C_JR,
		C_JALR,
		// RV64C
		C_ADDIW,
		C_SUBW,
		C_ADDW,
		C_LD,
		C_SD,
		C_LDSP,
		C_SDSP,
		// RV128C
		C_SRLI64,
		C_SRAI64,
		C_SLLI64,
		C_LQ,
		C_SQ,
		C_LQSP,
		C_SQSP,
		// RV32FC
		C_FLW,
		C_FSW,
		C_FLWSP,
		C_FSWSP,
		// RV32DC
		C_FLD,
		C_FSD,
		C_FLDSP,
		C_FSDSP,
		// RV32A
		LR_W,
		SC_W,
		AMOSWAP_W,
		AMOADD_W,
		AMOAND_W,
		AMOOR_W,
		AMOXOR_W,
		AMOMIN_W,
		AMOMAX_W,
		AMOMINU_W,
		AMOMAXU_W,
		// RV64A
		LR_D,
		SC_D,
		AMOSWAP_D,
		AMOADD_D,
		AMOAND_D,
		AMOOR_D,
		AMOXOR_D,
		AMOMIN_D,
		AMOMAX_D,
		AMOMINU_D,
		AMOMAXU_D,
		// Supervisor instruction
		DRET,
		MRET,
		URET,
		SRET,
		WFI,
		SFENCE_VMA,
		// You can add other instructions here
		INVALID_INSTR
	} riscv_instr_name_t;
	
	typedef enum bit [4:0] {
		ZERO = 5'b00000,
		RA,
		SP,
		GP,
		TP,
		T0,
		T1,
		T2,
		S0,
		S1,
		A0,
		A1,
		A2,
		A3,
		A4,
		A5,
		A6,
		A7,
		S2,
		S3,
		S4,
		S5,
		S6,
		S7,
		S8,
		S9,
		S10,
		S11,
		T3,
		T4,
		T5,
		T6
	} riscv_reg_t;

	typedef enum integer {
		J_FORMAT,
		U_FORMAT,
		I_FORMAT,
		I_FORMAT_SHIFT,
		B_FORMAT,
		R_FORMAT,
		S_FORMAT,
		CI_FORMAT,
		CB_FORMAT,
		CJ_FORMAT,
		CR_FORMAT,
		CL_FORMAT,
		CS_FORMAT,
		CSS_FORMAT,
		CIW_FORMAT
	} riscv_instr_format_t;

	typedef enum bit [3:0] {
		LOAD = 0,
		STORE,
		SHIFT,
		ARITHMETIC,
		LOGICAL,
		COMPARE,
		BRANCH,
		JUMP,
		SYNCH,
		SYSTEM,
		COUNTER,
		CSR,
		CHANGELEVEL,
		TRAP,
		INTERRUPT,
		AMO
	} riscv_instr_cateogry_t;
	
endpackage

`endif