function instruction_base_si sb_predictor::sb_calc_exp (instruction_base_si t);
	
	//instruction_base_si tr = instruction_base_si::type_id::create("tr");
	
	//`uvm_info(get_type_name(), t.convert2string(), UVM_HIGH)
	//tr.copy(t);

	//tr.address = 0;
	return(null);
endfunction 