function load_instruction_si sb_predictor::sb_calc_exp (load_instruction_si t);
	
	//load_instruction_si tr = load_instruction_si::type_id::create("tr");
	
	//`uvm_info(get_type_name(), t.convert2string(), UVM_HIGH)
	//tr.copy(t);

	//tr.address = 0;
	return(null);
endfunction 