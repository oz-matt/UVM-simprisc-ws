function arithmetic_instruction_si sb_predictor::sb_calc_exp (arithmetic_instruction_si t);
	
	//arithmetic_instruction_si tr = arithmetic_instruction_si::type_id::create("tr");
	
	//`uvm_info(get_type_name(), t.convert2string(), UVM_HIGH)
	//tr.copy(t);

	//tr.address = 0;
	return(null);
endfunction 