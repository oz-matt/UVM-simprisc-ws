`ifndef IGEN_UTILS
`define IGEN_UTILS

package igen_utils;
	
	`include "src/seq_items/asmutils.sv"
	
endpackage

`endif
